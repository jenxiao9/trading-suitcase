`ifndef BSH
`define BSH
parameter BSMODS = 1
parameter parameter DATASIZE = 224;
`endif